LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;
 
ENTITY Testbench_Data_Mem IS
END Testbench_Data_Mem;
 
ARCHITECTURE behavior OF Testbench_Data_Mem IS
 
-- Component Declaration for the Unit Under Test (UUT)

component Data_Mem
 port (Address: in STD_LOGIC_VECTOR (31 downto 0);
		 Write_Data: in STD_LOGIC_VECTOR (31 downto 0);
		 memWrite, memRead: in STD_LOGIC;
		 clk: in STD_LOGIC;
		 Read_Data: out STD_LOGIC_VECTOR (31 downto 0)); 
end component;
 
 constant Clock_Frequency: integer := 1e6; --1MHz
 constant Clock_Period: time := 1000 ms / Clock_Frequency;	--Clock Period is 1 us at 1MHz frequency
 
-- Inputs
 signal Address: STD_LOGIC_VECTOR (31 downto 0);
 signal Write_Data: STD_LOGIC_VECTOR (31 downto 0);
 signal memWrite, memRead: STD_LOGIC;
 signal CLK: STD_LOGIC := '0';
 
-- Outputs
 signal Read_Data: STD_LOGIC_VECTOR (31 downto 0); 
 
BEGIN
 
 -- Instantiate the Unit Under Test (UUT)
 uut: Data_Mem PORT MAP (
 Address => Address,
 Write_Data => Write_Data,
 memWrite => memWrite,
 memRead => memRead,
 clk => CLK,
 Read_Data => Read_Data
 );
 
 clk_process :process
   begin
		clk <= not clk;
		wait for Clock_Period/2;
  end process;
 
-- Stimulus process: no stimulus so runs through once
 stim_proc: process
 begin
 
 memWrite <= '1';
 
 Address <= std_logic_vector(to_unsigned(4, 32));
 Write_Data <= std_logic_vector(to_unsigned(333333333, 32));
 wait for Clock_Period;
 
 memWrite <= '1';
 
 Address <= std_logic_vector(to_unsigned(28, 32));
 Write_Data <= std_logic_vector(to_unsigned(555555555, 32));
 wait for Clock_Period;
 
 memWrite <= '0';
 
 Address <= std_logic_vector(to_unsigned(4, 32));
 Write_Data <= std_logic_vector(to_unsigned(11, 32));
 wait for Clock_Period;
 
 memRead <= '1'; 
 Address <= std_logic_vector(to_unsigned(28, 32));
 
 wait;
 end process;
 
END;
